`timescale 1ns/1ps

module poker(type, i0, i1, i2, i3, i4);
//DO NOT CHANGE!
	input  [5:0] i0, i1, i2, i3, i4;
	output [3:0] type;
//---------------------------------------------------
	EO en1(F40, i0[4], i1[4]);
	EO en2(F41, i1[4], i2[4]);
	EO en3(F42, i2[4], i3[4]);
	EO en4(F43, i3[4], i4[4]);
	OR4 fand1(F4, F40, F41, F42, F43);
	
	EO en5(F50, i0[5], i1[5]);
	EO en6(F51, i1[5], i2[5]);
	EO en7(F52, i2[5], i3[5]);
	EO en8(F53, i3[5], i4[5]);
	OR4 fand2(F5, F50, F51, F52, F53);

	NR2 fand3(FLOWER, F4, F5);
	IV FNAND3(NF, FLOWER);

	IV inv03(i03b, i0[3]);
	IV inv02(i02b, i0[2]);
	IV inv01(i01b, i0[1]);
	IV inv00(i00b, i0[0]);
	AN4 W013(Y013, i0[0], i01b, i0[2], i0[3]);
	AN4 W012(Y012, i00b, i01b, i0[2], i0[3]);
	AN4 W011(Y011, i0[0], i0[1], i02b, i0[3]);
	AN4 W010(Y010, i00b, i0[1], i02b, i0[3]);
	AN4 W09(Y09, i0[0], i01b, i02b, i0[3]);
	AN4 W08(Y08, i00b, i01b, i02b, i0[3]);
	AN4 W07(Y07, i0[0], i0[1], i0[2], i03b);
	AN4 W06(Y06, i00b, i0[1], i0[2], i03b);
	AN4 W05(Y05, i0[0], i01b, i0[2], i03b);
	AN4 W04(Y04, i00b, i01b, i0[2], i03b);
	AN4 W03(Y03, i0[0], i0[1], i02b, i03b);
	AN4 W02(Y02, i00b, i0[1], i02b, i03b);
	AN4 W01(Y01, i0[0], i01b, i02b, i03b);

	IV inv13(i13b, i1[3]);
	IV inv12(i12b, i1[2]);
	IV inv11(i11b, i1[1]);
	IV inv10(i10b, i1[0]);
	AN4 W113(Y113, i1[0], i11b, i1[2], i1[3]);
	AN4 W112(Y112, i10b, i11b, i1[2], i1[3]);
	AN4 W111(Y111, i1[0], i1[1], i12b, i1[3]);
	AN4 W110(Y110, i10b, i1[1], i12b, i1[3]);
	AN4 W19(Y19, i1[0], i11b, i12b, i1[3]);
	AN4 W18(Y18, i10b, i11b, i12b, i1[3]);
	AN4 W17(Y17, i1[0], i1[1], i1[2], i13b);
	AN4 W16(Y16, i10b, i1[1], i1[2], i13b);
	AN4 W15(Y15, i1[0], i11b, i1[2], i13b);
	AN4 W14(Y14, i10b, i11b, i1[2], i13b);
	AN4 W13(Y13, i1[0], i1[1], i12b, i13b);
	AN4 W12(Y12, i10b, i1[1], i12b, i13b);
	AN4 W11(Y11, i1[0], i11b, i12b, i13b);

	IV inv23(i23b, i2[3]);
	IV inv22(i22b, i2[2]);
	IV inv21(i21b, i2[1]);
	IV inv20(i20b, i2[0]);
	AN4 W213(Y213, i2[0], i21b, i2[2], i2[3]);
	AN4 W212(Y212, i20b, i21b, i2[2], i2[3]);
	AN4 W211(Y211, i2[0], i2[1], i22b, i2[3]);
	AN4 W210(Y210, i20b, i2[1], i22b, i2[3]);
	AN4 W29(Y29, i2[0], i21b, i22b, i2[3]);
	AN4 W28(Y28, i20b, i21b, i22b, i2[3]);
	AN4 W27(Y27, i2[0], i2[1], i2[2], i23b);
	AN4 W26(Y26, i20b, i2[1], i2[2], i23b);
	AN4 W25(Y25, i2[0], i21b, i2[2], i23b);
	AN4 W24(Y24, i20b, i21b, i2[2], i23b);
	AN4 W23(Y23, i2[0], i2[1], i22b, i23b);
	AN4 W22(Y22, i20b, i2[1], i22b, i23b);
	AN4 W21(Y21, i2[0], i21b, i22b, i23b);

	IV inv33(i33b, i3[3]);
	IV inv32(i32b, i3[2]);
	IV inv31(i31b, i3[1]);
	IV inv30(i30b, i3[0]);
	AN4 W313(Y313, i3[0], i31b, i3[2], i3[3]);
	AN4 W312(Y312, i30b, i31b, i3[2], i3[3]);
	AN4 W311(Y311, i3[0], i3[1], i32b, i3[3]);
	AN4 W310(Y310, i30b, i3[1], i32b, i3[3]);
	AN4 W39(Y39, i3[0], i31b, i32b, i3[3]);
	AN4 W38(Y38, i30b, i31b, i32b, i3[3]);
	AN4 W37(Y37, i3[0], i3[1], i3[2], i33b);
	AN4 W36(Y36, i30b, i3[1], i3[2], i33b);
	AN4 W35(Y35, i3[0], i31b, i3[2], i33b);
	AN4 W34(Y34, i30b, i31b, i3[2], i33b);
	AN4 W33(Y33, i3[0], i3[1], i32b, i33b);
	AN4 W32(Y32, i30b, i3[1], i32b, i33b);
	AN4 W31(Y31, i3[0], i31b, i32b, i33b);

	IV inv43(i43b, i4[3]);
	IV inv42(i42b, i4[2]);
	IV inv41(i41b, i4[1]);
	IV inv40(i40b, i4[0]);
	AN4 W413(Y413, i4[0], i41b, i4[2], i4[3]);
	AN4 W412(Y412, i40b, i41b, i4[2], i4[3]);
	AN4 W411(Y411, i4[0], i4[1], i42b, i4[3]);
	AN4 W410(Y410, i40b, i4[1], i42b, i4[3]);
	AN4 W49(Y49, i4[0], i41b, i42b, i4[3]);
	AN4 W48(Y48, i40b, i41b, i42b, i4[3]);
	AN4 W47(Y47, i4[0], i4[1], i4[2], i43b);
	AN4 W46(Y46, i40b, i4[1], i4[2], i43b);
	AN4 W45(Y45, i4[0], i41b, i4[2], i43b);
	AN4 W44(Y44, i40b, i41b, i4[2], i43b);
	AN4 W43(Y43, i4[0], i4[1], i42b, i43b);
	AN4 W42(Y42, i40b, i4[1], i42b, i43b);
	AN4 W41(Y41, i4[0], i41b, i42b, i43b);

	OR3 Yo130(YOR130, Y013, Y113, Y213);
	OR3 Yo131(YOR131, YOR130, Y313, Y413);
	OR3 Yo120(YOR120, Y012, Y112, Y212);
	OR3 Yo121(YOR121, YOR120, Y312, Y412);
	OR3 Yo110(YOR110, Y011, Y111, Y211);
	OR3 Yo111(YOR111, YOR110, Y311, Y411);
	OR3 Yo100(YOR100, Y010, Y110, Y210);
	OR3 Yo101(YOR101, YOR100, Y310, Y410);
	OR3 Yo90(YOR90, Y09, Y19, Y29);
	OR3 Yo91(YOR91, YOR90, Y39, Y49);
	OR3 Yo80(YOR80, Y08, Y18, Y28);
	OR3 Yo81(YOR81, YOR80, Y38, Y48);
	OR3 Yo70(YOR70, Y07, Y17, Y27);
	OR3 Yo71(YOR71, YOR70, Y37, Y47);
	OR3 Yo60(YOR60, Y06, Y16, Y26);
	OR3 Yo61(YOR61, YOR60, Y36, Y46);
	OR3 Yo50(YOR50, Y05, Y15, Y25);
	OR3 Yo51(YOR51, YOR50, Y35, Y45);
	OR3 Yo40(YOR40, Y04, Y14, Y24);
	OR3 Yo41(YOR41, YOR40, Y34, Y44);
	OR3 Yo30(YOR30, Y03, Y13, Y23);
	OR3 Yo31(YOR31, YOR30, Y33, Y43);
	OR3 Yo20(YOR20, Y02, Y12, Y22);
	OR3 Yo21(YOR21, YOR20, Y32, Y42);
	OR3 Yo10(YOR10, Y01, Y11, Y21);
	OR3 Yo11(YOR11, YOR10, Y31, Y41);

	AN3 AKB140(H14, YOR11, YOR131, YOR121);
	AN3 AKB141(G14, H14, YOR111, YOR101);
	AN3 AKB130(H13, YOR131, YOR121, YOR111);
	AN3 AKB131(G13, H13, YOR101, YOR91);
	AN3 AKB120(H12, YOR121, YOR111, YOR101);
	AN3 AKB121(G12, H12, YOR91, YOR81);
	AN3 AKB110(H11, YOR111, YOR101, YOR91);
	AN3 AKB111(G11, H11, YOR81, YOR71);
	AN3 AKB100(H10, YOR101, YOR91, YOR81);
	AN3 AKB101(G10, H10, YOR71, YOR61);
	AN3 AKB90(H9, YOR91, YOR81, YOR71);
	AN3 AKB91(G9, H9, YOR61, YOR51);
	AN3 AKB80(H8, YOR81, YOR71, YOR61);
	AN3 AKB81(G8, H8, YOR51, YOR41);
	AN3 AKB70(H7, YOR71, YOR61, YOR51);
	AN3 AKB71(G7, H7, YOR41, YOR31);
	AN3 AKB60(H6, YOR61, YOR51, YOR41);
	AN3 AKB61(G6, H6, YOR31, YOR21);
	AN3 AKB50(H5, YOR51, YOR41, YOR31);
	AN3 AKB51(G5, H5, YOR21, YOR11);

	NR3 KC0(CH1, G13, G12, G11);
	NR3 KC1(CH2, G10, G9, G8);
	NR3 KC2(CH3, G7, G6, G5);
	IV KKG(NG14, G14);
	ND4 KC(CHILL, NG14, CH1, CH2, CH3);

	HA1 HA130(C113, S013, Y013, Y113);
	FA1 FA130(C413, S313, Y213, Y313, Y413);
	HA1 HA131(C213, A130, S313, S013);
	FA1 FA131(A132, A131, C213, C113, C413);
	HA1 HA120(C112, S012, Y012, Y112);
	FA1 FA120(C412, S312, Y212, Y312, Y412);
	HA1 HA121(C212, A120, S312, S012);
	FA1 FA121(A122, A121, C212, C112, C412);
	HA1 HA110(C111, S011, Y011, Y111);
	FA1 FA110(C411, S311, Y211, Y311, Y411);
	HA1 HA111(C211, A110, S311, S011);
	FA1 FA111(A112, A111, C211, C111, C411);
	HA1 HA100(C110, S010, Y010, Y110);
	FA1 FA100(C410, S310, Y210, Y310, Y410);
	HA1 HA101(C210, A100, S310, S010);
	FA1 FA101(A102, A101, C210, C110, C410);
	HA1 HA90(C19, S09, Y09, Y19);
	FA1 FA90(C49, S39, Y29, Y39, Y49);
	HA1 HA91(C29, A90, S39, S09);
	FA1 FA91(A92, A91, C29, C19, C49);
	HA1 HA80(C18, S08, Y08, Y18);
	FA1 FA80(C48, S38, Y28, Y38, Y48);
	HA1 HA81(C28, A80, S38, S08);
	FA1 FA81(A82, A81, C28, C18, C48);
	HA1 HA70(C17, S07, Y07, Y17);
	FA1 FA70(C47, S37, Y27, Y37, Y47);
	HA1 HA71(C27, A70, S37, S07);
	FA1 FA71(A72, A71, C27, C17, C47);
	HA1 HA60(C16, S06, Y06, Y16);
	FA1 FA60(C46, S36, Y26, Y36, Y46);
	HA1 HA61(C26, A60, S36, S06);
	FA1 FA61(A62, A61, C26, C16, C46);
	HA1 HA50(C15, S05, Y05, Y15);
	FA1 FA50(C45, S35, Y25, Y35, Y45);
	HA1 HA51(C25, A50, S35, S05);
	FA1 FA51(A52, A51, C25, C15, C45);
	HA1 HA40(C14, S04, Y04, Y14);
	FA1 FA40(C44, S34, Y24, Y34, Y44);
	HA1 HA41(C24, A40, S34, S04);
	FA1 FA41(A42, A41, C24, C14, C44);
	HA1 HA30(C13, S03, Y03, Y13);
	FA1 FA30(C43, S33, Y23, Y33, Y43);
	HA1 HA31(C23, A30, S33, S03);
	FA1 FA31(A32, A31, C23, C13, C43);
	HA1 HA20(C12, S02, Y02, Y12);
	FA1 FA20(C42, S32, Y22, Y32, Y42);
	HA1 HA21(C22, A20, S32, S02);
	FA1 FA21(A22, A21, C22, C12, C42);
	HA1 HA10(C11, S01, Y01, Y11);
	FA1 FA10(C41, S31, Y21, Y31, Y41);
	HA1 HA11(C21, A10, S31, S01);
	FA1 FA11(A12, A11, C21, C11, C41);

	ND2 KAND13(K13, A130, A131);
	ND2 KAND12(K12, A120, A121);
	ND2 KAND11(K11, A110, A111);
	ND2 KAND10(K10, A100, A101);
	ND2 KAND9(K9, A90, A91);
	ND2 KAND8(K8, A80, A81);
	ND2 KAND7(K7, A70, A71);
	ND2 KAND6(K6, A60, A61);
	ND2 KAND5(K5, A50, A51);
	ND2 KAND4(K4, A40, A41);
	ND2 KAND3(K3, A30, A31);
	ND2 KAND2(K2, A20, A21);
	AN2 KAND1(K1, A10, A11);
	ND4 KKOR0(KK1, K13, K12, K11, K10);
	ND4 KKOR1(KK2, K9, K8, K7, K6);
	ND4 KKOR2(KK3, K5, K4, K3, K2);
	OR4 KKOR(ANBN, KK1, KK2, KK3, K1);
	
	//EO3 KXOR12(KX12, A131, A121, A111);
	EO FG121(FFG1, A131, A121);
	EO FG122(KX12, FFG1, A111);
	//EO3 KXOR8(KX8, A101, A91, A81);
	EO FG81(FFG2, A101, A91);
	EO FG82(KX8, FFG2, A81);
	//EO3 KXOR5(KX5, A71, A61, A51);
	EO FG51(FFG3, A71, A61);
	EO FG52(KX5, FFG3, A51);
	//EO3 KXOR2(KX2, A41, A31, A21);
	EO FG21(FFG4, A41, A31);
	EO FG22(KX2, FFG4, A21);
	//EO3 KXOR1(BNXOR, KX2, A11, KX0);
	EO FG11(FFG5, KX2, A11);
	EO FG12(BNXOR, FFG5, KX0);
	EO3 KKXOR0(KX0, KX12, KX8, KX5);
	EO FG1(FFG01, KX12, KX8);
	EO FG2(KX0, FFG01, KX5);
	IV LA3(NBNXOR, BNXOR);

	OR4 KOR10(B0, A131, A121, A111, A101);
	OR4 KOR6(B1, A91, A81, A71, A61);
	OR4 KOR2(B2, A51, A41, A31, A21);
	OR4 KOR(BNOR, B0, B1, B2, A11);

	OR4 COR0(C1, A132, A122, A112, A102);
	OR4 COR1(C2, A92, A82, A72, A62);
	OR4 COR2(C3, A52, A42, A32, A22);
	OR4 COR(CNOR, C1, C2, C3, A12);

	AN2 TT1(T1, FLOWER, NCHILL);
	IV IVANBN(NANBN, ANBN);
	IV IVBNOR(NBNOR, BNOR);
	ND2 QAN1(Q41, NBNXOR, CNOR);
	ND2 QAN2(Q32, ANBN, NBNXOR);
	ND2 QAN3(Q311, ANBN, BNXOR);
	ND2 QAN4(Q221, NBNXOR, BNOR);
	ND2 QAN5(Q2111, NANBN, BNXOR);
	ND2 QAN6(Q11111, NBNOR, T1);
	IV IVC(NCHILL, CHILL);
	AN2 QAN7(type[3], CHILL, FLOWER);
	ND2 QAN8(J0, NF, CHILL);
	ND4 ANS2(type[2], Q11111, Q41, Q32, J0);
	ND4 ANS1(type[1], Q41, Q32, Q311, Q221);
	ND4 ANS0(type[0], Q41, Q311, Q2111, Q11111);

endmodule