`timescale 1ns/1ps

module poker(type, i0, i1, i2, i3, i4);
//DO NOT CHANGE!
	input  [5:0] i0, i1, i2, i3, i4;
	output [3:0] type;
//---------------------------------------------------
	EO en1(F40, i0[4], i1[4]);
	EO en2(F41, i1[4], i2[4]);
	EO en3(F42, i2[4], i3[4]);
	EO en4(F43, i3[4], i4[4]);
	OR4 fand1(F4, F40, F41, F42, F43);
	
	EO en5(F50, i0[5], i1[5]);
	EO en6(F51, i1[5], i2[5]);
	EO en7(F52, i2[5], i3[5]);
	EO en8(F53, i3[5], i4[5]);
	OR4 fand2(F5, F50, F51, F52, F53);

	NR2 fand3(FLOWER, F4, F5);
	IV FNAND3(NF, FLOWER);

	IV inv03(i03b, i0[3]);
	IV inv02(i02b, i0[2]);
	IV inv01(i01b, i0[1]);
	IV inv00(i00b, i0[0]);
	AN4 W013(Y013, i0[0], i01b, i0[2], i0[3]);
	AN4 W012(Y012, i00b, i01b, i0[2], i0[3]);
	AN4 W011(Y011, i0[0], i0[1], i02b, i0[3]);
	AN4 W010(Y010, i00b, i0[1], i02b, i0[3]);
	AN4 W09(Y09, i0[0], i01b, i02b, i0[3]);
	AN4 W08(Y08, i00b, i01b, i02b, i0[3]);
	AN4 W07(Y07, i0[0], i0[1], i0[2], i03b);
	AN4 W06(Y06, i00b, i0[1], i0[2], i03b);
	AN4 W05(Y05, i0[0], i01b, i0[2], i03b);
	AN4 W04(Y04, i00b, i01b, i0[2], i03b);
	AN4 W03(Y03, i0[0], i0[1], i02b, i03b);
	AN4 W02(Y02, i00b, i0[1], i02b, i03b);
	AN4 W01(Y01, i0[0], i01b, i02b, i03b);

	IV inv13(i13b, i1[3]);
	IV inv12(i12b, i1[2]);
	IV inv11(i11b, i1[1]);
	IV inv10(i10b, i1[0]);
	AN4 W113(Y113, i1[0], i11b, i1[2], i1[3]);
	AN4 W112(Y112, i10b, i11b, i1[2], i1[3]);
	AN4 W111(Y111, i1[0], i1[1], i12b, i1[3]);
	AN4 W110(Y110, i10b, i1[1], i12b, i1[3]);
	AN4 W19(Y19, i1[0], i11b, i12b, i1[3]);
	AN4 W18(Y18, i10b, i11b, i12b, i1[3]);
	AN4 W17(Y17, i1[0], i1[1], i1[2], i13b);
	AN4 W16(Y16, i10b, i1[1], i1[2], i13b);
	AN4 W15(Y15, i1[0], i11b, i1[2], i13b);
	AN4 W14(Y14, i10b, i11b, i1[2], i13b);
	AN4 W13(Y13, i1[0], i1[1], i12b, i13b);
	AN4 W12(Y12, i10b, i1[1], i12b, i13b);
	AN4 W11(Y11, i1[0], i11b, i12b, i13b);

	IV inv23(i23b, i2[3]);
	IV inv22(i22b, i2[2]);
	IV inv21(i21b, i2[1]);
	IV inv20(i20b, i2[0]);
	AN4 W213(Y213, i2[0], i21b, i2[2], i2[3]);
	AN4 W212(Y212, i20b, i21b, i2[2], i2[3]);
	AN4 W211(Y211, i2[0], i2[1], i22b, i2[3]);
	AN4 W210(Y210, i20b, i2[1], i22b, i2[3]);
	AN4 W29(Y29, i2[0], i21b, i22b, i2[3]);
	AN4 W28(Y28, i20b, i21b, i22b, i2[3]);
	AN4 W27(Y27, i2[0], i2[1], i2[2], i23b);
	AN4 W26(Y26, i20b, i2[1], i2[2], i23b);
	AN4 W25(Y25, i2[0], i21b, i2[2], i23b);
	AN4 W24(Y24, i20b, i21b, i2[2], i23b);
	AN4 W23(Y23, i2[0], i2[1], i22b, i23b);
	AN4 W22(Y22, i20b, i2[1], i22b, i23b);
	AN4 W21(Y21, i2[0], i21b, i22b, i23b);

	IV inv33(i33b, i3[3]);
	IV inv32(i32b, i3[2]);
	IV inv31(i31b, i3[1]);
	IV inv30(i30b, i3[0]);
	AN4 W313(Y313, i3[0], i31b, i3[2], i3[3]);
	AN4 W312(Y312, i30b, i31b, i3[2], i3[3]);
	AN4 W311(Y311, i3[0], i3[1], i32b, i3[3]);
	AN4 W310(Y310, i30b, i3[1], i32b, i3[3]);
	AN4 W39(Y39, i3[0], i31b, i32b, i3[3]);
	AN4 W38(Y38, i30b, i31b, i32b, i3[3]);
	AN4 W37(Y37, i3[0], i3[1], i3[2], i33b);
	AN4 W36(Y36, i30b, i3[1], i3[2], i33b);
	AN4 W35(Y35, i3[0], i31b, i3[2], i33b);
	AN4 W34(Y34, i30b, i31b, i3[2], i33b);
	AN4 W33(Y33, i3[0], i3[1], i32b, i33b);
	AN4 W32(Y32, i30b, i3[1], i32b, i33b);
	AN4 W31(Y31, i3[0], i31b, i32b, i33b);

	IV inv43(i43b, i4[3]);
	IV inv42(i42b, i4[2]);
	IV inv41(i41b, i4[1]);
	IV inv40(i40b, i4[0]);
	AN4 W413(Y413, i4[0], i41b, i4[2], i4[3]);
	AN4 W412(Y412, i40b, i41b, i4[2], i4[3]);
	AN4 W411(Y411, i4[0], i4[1], i42b, i4[3]);
	AN4 W410(Y410, i40b, i4[1], i42b, i4[3]);
	AN4 W49(Y49, i4[0], i41b, i42b, i4[3]);
	AN4 W48(Y48, i40b, i41b, i42b, i4[3]);
	AN4 W47(Y47, i4[0], i4[1], i4[2], i43b);
	AN4 W46(Y46, i40b, i4[1], i4[2], i43b);
	AN4 W45(Y45, i4[0], i41b, i4[2], i43b);
	AN4 W44(Y44, i40b, i41b, i4[2], i43b);
	AN4 W43(Y43, i4[0], i4[1], i42b, i43b);
	AN4 W42(Y42, i40b, i4[1], i42b, i43b);
	AN4 W41(Y41, i4[0], i41b, i42b, i43b);

	OR3 Yo130(YOR130, Y013, Y113, Y213);
	OR3 Yo131(YOR131, YOR130, Y313, Y413);
	OR3 Yo120(YOR120, Y012, Y112, Y212);
	OR3 Yo121(YOR121, YOR120, Y312, Y412);
	OR3 Yo110(YOR110, Y011, Y111, Y211);
	OR3 Yo111(YOR111, YOR110, Y311, Y411);
	OR3 Yo100(YOR100, Y010, Y110, Y210);
	OR3 Yo101(YOR101, YOR100, Y310, Y410);
	OR3 Yo90(YOR90, Y09, Y19, Y29);
	OR3 Yo91(YOR91, YOR90, Y39, Y49);
	OR3 Yo80(YOR80, Y08, Y18, Y28);
	OR3 Yo81(YOR81, YOR80, Y38, Y48);
	OR3 Yo70(YOR70, Y07, Y17, Y27);
	OR3 Yo71(YOR71, YOR70, Y37, Y47);
	OR3 Yo60(YOR60, Y06, Y16, Y26);
	OR3 Yo61(YOR61, YOR60, Y36, Y46);
	OR3 Yo50(YOR50, Y05, Y15, Y25);
	OR3 Yo51(YOR51, YOR50, Y35, Y45);
	OR3 Yo40(YOR40, Y04, Y14, Y24);
	OR3 Yo41(YOR41, YOR40, Y34, Y44);
	OR3 Yo30(YOR30, Y03, Y13, Y23);
	OR3 Yo31(YOR31, YOR30, Y33, Y43);
	OR3 Yo20(YOR20, Y02, Y12, Y22);
	OR3 Yo21(YOR21, YOR20, Y32, Y42);
	OR3 Yo10(YOR10, Y01, Y11, Y21);
	OR3 Yo11(YOR11, YOR10, Y31, Y41);

	AN3 AKB140(H14, YOR11, YOR131, YOR121);
	AN3 AKB141(G14, H14, YOR111, YOR101);
	AN3 AKB130(H13, YOR131, YOR121, YOR111);
	AN3 AKB131(G13, H13, YOR101, YOR91);
	AN3 AKB120(H12, YOR121, YOR111, YOR101);
	AN3 AKB121(G12, H12, YOR91, YOR81);
	AN3 AKB110(H11, YOR111, YOR101, YOR91);
	AN3 AKB111(G11, H11, YOR81, YOR71);
	AN3 AKB100(H10, YOR101, YOR91, YOR81);
	AN3 AKB101(G10, H10, YOR71, YOR61);
	AN3 AKB90(H9, YOR91, YOR81, YOR71);
	AN3 AKB91(G9, H9, YOR61, YOR51);
	AN3 AKB80(H8, YOR81, YOR71, YOR61);
	AN3 AKB81(G8, H8, YOR51, YOR41);
	AN3 AKB70(H7, YOR71, YOR61, YOR51);
	AN3 AKB71(G7, H7, YOR41, YOR31);
	AN3 AKB60(H6, YOR61, YOR51, YOR41);
	AN3 AKB61(G6, H6, YOR31, YOR21);
	AN3 AKB50(H5, YOR51, YOR41, YOR31);
	AN3 AKB51(G5, H5, YOR21, YOR11);

	NR3 KC0(CH1, G13, G12, G11);
	NR3 KC1(CH2, G10, G9, G8);
	NR3 KC2(CH3, G7, G6, G5);
	IV KKG(NG14, G14);
	ND4 KC(CHILL, NG14, CH1, CH2, CH3);

	ND3 PPA11(PA11, Y01, Y11, Y21);
	ND3 PPA12(PA12, Y11, Y21, Y31);
	ND3 PPA13(PA13, Y21, Y31, Y41);
	ND3 PPA14(PA14, Y11, Y31, Y41);
	ND3 PPA15(PA15, Y11, Y21, Y41);
	ND3 PPA16(PA16, Y01, Y31, Y41);
	ND3 PPA17(PA17, Y01, Y21, Y41);
	ND3 PPA18(PA18, Y01, Y21, Y31);
	ND3 PPA19(PA19, Y01, Y11, Y41);
	ND3 PPA110(PA110, Y01, Y11, Y31);
	AN4 PPO11(PO11, PA11, PA12, PA13, PA14);
	AN4 PPO12(PO12, PA15, PA16, PA17, PA18);
	ND4 PPO13(PO13, PA19, PA110, PO11, PO12);
	
	ND3 PPA21(PA21, Y02, Y12, Y22);
	ND3 PPA22(PA22, Y12, Y22, Y32);
	ND3 PPA23(PA23, Y22, Y32, Y42);
	ND3 PPA24(PA24, Y12, Y32, Y42);
	ND3 PPA25(PA25, Y12, Y22, Y42);
	ND3 PPA26(PA26, Y02, Y32, Y42);
	ND3 PPA27(PA27, Y02, Y22, Y42);
	ND3 PPA28(PA28, Y02, Y22, Y32);
	ND3 PPA29(PA29, Y02, Y12, Y42);
	ND3 PPA210(PA210, Y02, Y12, Y32);
	AN4 PPO21(PO21, PA21, PA22, PA23, PA24);
	AN4 PPO22(PO22, PA25, PA26, PA27, PA28);
	ND4 PPO23(PO23, PA29, PA210, PO21, PO22);

	ND3 PPA31(PA31, Y03, Y13, Y23);
	ND3 PPA32(PA32, Y13, Y23, Y33);
	ND3 PPA33(PA33, Y23, Y33, Y43);
	ND3 PPA34(PA34, Y13, Y33, Y43);
	ND3 PPA35(PA35, Y13, Y23, Y43);
	ND3 PPA36(PA36, Y03, Y33, Y43);
	ND3 PPA37(PA37, Y03, Y23, Y43);
	ND3 PPA38(PA38, Y03, Y23, Y33);
	ND3 PPA39(PA39, Y03, Y13, Y43);
	ND3 PPA310(PA310, Y03, Y13, Y33);
	AN4 PPO31(PO31, PA31, PA32, PA33, PA34);
	AN4 PPO32(PO32, PA35, PA36, PA37, PA38);
	ND4 PPO33(PO33, PA39, PA310, PO31, PO32);

	ND3 PPA41(PA41, Y04, Y14, Y24);
	ND3 PPA42(PA42, Y14, Y24, Y34);
	ND3 PPA43(PA43, Y24, Y34, Y44);
	ND3 PPA44(PA44, Y14, Y34, Y44);
	ND3 PPA45(PA45, Y14, Y24, Y44);
	ND3 PPA46(PA46, Y04, Y34, Y44);
	ND3 PPA47(PA47, Y04, Y24, Y44);
	ND3 PPA48(PA48, Y04, Y24, Y34);
	ND3 PPA49(PA49, Y04, Y14, Y44);
	ND3 PPA410(PA410, Y04, Y14, Y34);
	AN4 PPO41(PO41, PA41, PA42, PA43, PA44);
	AN4 PPO42(PO42, PA45, PA46, PA47, PA48);
	ND4 PPO43(PO43, PA49, PA410, PO41, PO42);

	ND3 PPA51(PA51, Y05, Y15, Y25);
	ND3 PPA52(PA52, Y15, Y25, Y35);
	ND3 PPA53(PA53, Y25, Y35, Y45);
	ND3 PPA54(PA54, Y15, Y35, Y45);
	ND3 PPA55(PA55, Y15, Y25, Y45);
	ND3 PPA56(PA56, Y05, Y35, Y45);
	ND3 PPA57(PA57, Y05, Y25, Y45);
	ND3 PPA58(PA58, Y05, Y25, Y35);
	ND3 PPA59(PA59, Y05, Y15, Y45);
	ND3 PPA510(PA510, Y05, Y15, Y35);
	AN4 PPO51(PO51, PA51, PA52, PA53, PA54);
	AN4 PPO52(PO52, PA55, PA56, PA57, PA58);
	ND4 PPO53(PO53, PA59, PA510, PO51, PO52);

	ND3 PPA61(PA61, Y06, Y16, Y26);
	ND3 PPA62(PA62, Y16, Y26, Y36);
	ND3 PPA63(PA63, Y26, Y36, Y46);
	ND3 PPA64(PA64, Y16, Y36, Y46);
	ND3 PPA65(PA65, Y16, Y26, Y46);
	ND3 PPA66(PA66, Y06, Y36, Y46);
	ND3 PPA67(PA67, Y06, Y26, Y46);
	ND3 PPA68(PA68, Y06, Y26, Y36);
	ND3 PPA69(PA69, Y06, Y16, Y46);
	ND3 PPA610(PA610, Y06, Y16, Y36);
	AN4 PPO61(PO61, PA61, PA62, PA63, PA64);
	AN4 PPO62(PO62, PA65, PA66, PA67, PA68);
	ND4 PPO63(PO63, PA69, PA610, PO61, PO62);

	ND3 PPA71(PA71, Y07, Y17, Y27);
	ND3 PPA72(PA72, Y17, Y27, Y37);
	ND3 PPA73(PA73, Y27, Y37, Y47);
	ND3 PPA74(PA74, Y17, Y37, Y47);
	ND3 PPA75(PA75, Y17, Y27, Y47);
	ND3 PPA76(PA76, Y07, Y37, Y47);
	ND3 PPA77(PA77, Y07, Y27, Y47);
	ND3 PPA78(PA78, Y07, Y27, Y37);
	ND3 PPA79(PA79, Y07, Y17, Y47);
	ND3 PPA710(PA710, Y07, Y17, Y37);
	AN4 PPO71(PO71, PA71, PA72, PA73, PA74);
	AN4 PPO72(PO72, PA75, PA76, PA77, PA78);
	ND4 PPO73(PO73, PA79, PA710, PO71, PO72);

	ND3 PPA81(PA81, Y08, Y18, Y28);
	ND3 PPA82(PA82, Y18, Y28, Y38);
	ND3 PPA83(PA83, Y28, Y38, Y48);
	ND3 PPA84(PA84, Y18, Y38, Y48);
	ND3 PPA85(PA85, Y18, Y28, Y48);
	ND3 PPA86(PA86, Y08, Y38, Y48);
	ND3 PPA87(PA87, Y08, Y28, Y48);
	ND3 PPA88(PA88, Y08, Y28, Y38);
	ND3 PPA89(PA89, Y08, Y18, Y48);
	ND3 PPA810(PA810, Y08, Y18, Y38);
	AN4 PPO81(PO81, PA81, PA82, PA83, PA84);
	AN4 PPO82(PO82, PA85, PA86, PA87, PA88);
	ND4 PPO83(PO83, PA89, PA810, PO81, PO82);

	ND3 PPA91(PA91, Y09, Y19, Y29);
	ND3 PPA92(PA92, Y19, Y29, Y39);
	ND3 PPA93(PA93, Y29, Y39, Y49);
	ND3 PPA94(PA94, Y19, Y39, Y49);
	ND3 PPA95(PA95, Y19, Y29, Y49);
	ND3 PPA96(PA96, Y09, Y39, Y49);
	ND3 PPA97(PA97, Y09, Y29, Y49);
	ND3 PPA98(PA98, Y09, Y29, Y39);
	ND3 PPA99(PA99, Y09, Y19, Y49);
	ND3 PPA910(PA910, Y09, Y19, Y39);
	AN4 PPO91(PO91, PA91, PA92, PA93, PA94);
	AN4 PPO92(PO92, PA95, PA96, PA97, PA98);
	ND4 PPO93(PO93, PA99, PA910, PO91, PO92);

	ND3 PPA101(PA101, Y010, Y110, Y210);
	ND3 PPA102(PA102, Y110, Y210, Y310);
	ND3 PPA103(PA103, Y210, Y310, Y410);
	ND3 PPA104(PA104, Y110, Y310, Y410);
	ND3 PPA105(PA105, Y110, Y210, Y410);
	ND3 PPA106(PA106, Y010, Y310, Y410);
	ND3 PPA107(PA107, Y010, Y210, Y410);
	ND3 PPA108(PA108, Y010, Y210, Y310);
	ND3 PPA109(PA109, Y010, Y110, Y410);
	ND3 PPA1010(PA1010, Y010, Y110, Y310);
	AN4 PPO101(PO101, PA101, PA102, PA103, PA104);
	AN4 PPO102(PO102, PA105, PA106, PA107, PA108);
	ND4 PPO103(PO103, PA109, PA1010, PO101, PO102);

	AN3 PPA111(PA111, Y011, Y111, Y211);
	AN3 PPA112(PA112, Y111, Y211, Y311);
	AN3 PPA113(PA113, Y211, Y311, Y411);
	AN3 PPA114(PA114, Y111, Y311, Y411);
	AN3 PPA115(PA115, Y111, Y211, Y411);
	AN3 PPA116(PA116, Y011, Y311, Y411);
	AN3 PPA117(PA117, Y011, Y211, Y411);
	AN3 PPA118(PA118, Y011, Y211, Y311);
	AN3 PPA119(PA119, Y011, Y111, Y411);
	AN3 PPA1110(PA1110, Y011, Y111, Y311);
	OR4 PPO111(PO111, PA111, PA112, PA113, PA114);
	OR4 PPO112(PO112, PA115, PA116, PA117, PA118);
	OR4 PPO113(PO113, PA119, PA1110, PO111, PO112);

	ND3 PPA121(PA121, Y012, Y112, Y212);
	ND3 PPA122(PA122, Y112, Y212, Y312);
	ND3 PPA123(PA123, Y212, Y312, Y412);
	ND3 PPA124(PA124, Y112, Y312, Y412);
	ND3 PPA125(PA125, Y112, Y212, Y412);
	ND3 PPA126(PA126, Y012, Y312, Y412);
	ND3 PPA127(PA127, Y012, Y212, Y412);
	ND3 PPA128(PA128, Y012, Y212, Y312);
	ND3 PPA129(PA129, Y012, Y112, Y412);
	ND3 PPA1210(PA1210, Y012, Y112, Y312);
	AN4 PPO121(PO121, PA121, PA122, PA123, PA124);
	AN4 PPO122(PO122, PA125, PA126, PA127, PA128);
	ND4 PPO123(PO123, PA129, PA1210, PO121, PO122);

	ND3 PPA131(PA131, Y013, Y113, Y213);
	ND3 PPA132(PA132, Y113, Y213, Y313);
	ND3 PPA133(PA133, Y213, Y313, Y413);
	ND3 PPA134(PA134, Y113, Y313, Y413);
	ND3 PPA135(PA135, Y113, Y213, Y413);
	ND3 PPA136(PA136, Y013, Y313, Y413);
	ND3 PPA137(PA137, Y013, Y213, Y413);
	ND3 PPA138(PA138, Y013, Y213, Y313);
	ND3 PPA139(PA139, Y013, Y113, Y413);
	ND3 PPA1310(PA1310, Y013, Y113, Y313);
	AN4 PPO131(PO131, PA131, PA132, PA133, PA134);
	AN4 PPO132(PO132, PA135, PA136, PA137, PA138);
	ND4 PPO133(PO133, PA139, PA1310, PO131, PO132);

	NR3 PPS11(PS11, PO13, PO23, PO33);
	NR3 PPS21(PS21, PO43, PO53, PO63);
	NR3 PPS31(PS31, PO73, PO83, PO93);
	NR4 PPS41(PS41, PO103, PO113, PO123, PO133);
	ND4 PPS51(Q3, PS11, PS21, PS31, PS41);
	AN4 PPS511(NQ3, PS11, PS21, PS31, PS41);

	ND2 PPAA11(PAA11, Y01, Y11);
	ND2 PPAA12(PAA12, Y01, Y21);
	ND2 PPAA13(PAA13, Y01, Y31);
	ND2 PPAA14(PAA14, Y01, Y41);
	ND2 PPAA15(PAA15, Y11, Y21);
	ND2 PPAA16(PAA16, Y11, Y31);
	ND2 PPAA17(PAA17, Y11, Y41);
	ND2 PPAA18(PAA18, Y21, Y31);
	ND2 PPAA19(PAA19, Y21, Y41);
	ND2 PPAA110(PAA110, Y31, Y41);
	AN4 PPOO11(POO11, PAA11, PAA12, PAA13, PAA14);
	AN4 PPOO12(POO12, PAA15, PAA16, PAA17, PAA18);
	ND4 PPOO13(POO13, PAA19, PAA110, POO11, POO12);

	ND2 PPAA21(PAA21, Y02, Y12);
	ND2 PPAA22(PAA22, Y02, Y22);
	ND2 PPAA23(PAA23, Y02, Y32);
	ND2 PPAA24(PAA24, Y02, Y42);
	ND2 PPAA25(PAA25, Y12, Y22);
	ND2 PPAA26(PAA26, Y12, Y32);
	ND2 PPAA27(PAA27, Y12, Y42);
	ND2 PPAA28(PAA28, Y22, Y32);
	ND2 PPAA29(PAA29, Y22, Y42);
	ND2 PPAA210(PAA210, Y32, Y42);
	AN4 PPOO21(POO21, PAA21, PAA22, PAA23, PAA24);
	AN4 PPOO22(POO22, PAA25, PAA26, PAA27, PAA28);
	ND4 PPOO23(POO23, PAA29, PAA210, POO21, POO22);

	ND2 PPAA31(PAA31, Y03, Y13);
	ND2 PPAA32(PAA32, Y03, Y23);
	ND2 PPAA33(PAA33, Y03, Y33);
	ND2 PPAA34(PAA34, Y03, Y43);
	ND2 PPAA35(PAA35, Y13, Y23);
	ND2 PPAA36(PAA36, Y13, Y33);
	ND2 PPAA37(PAA37, Y13, Y43);
	ND2 PPAA38(PAA38, Y23, Y33);
	ND2 PPAA39(PAA39, Y23, Y43);
	ND2 PPAA310(PAA310, Y33, Y43);
	AN4 PPOO31(POO31, PAA31, PAA32, PAA33, PAA34);
	AN4 PPOO32(POO32, PAA35, PAA36, PAA37, PAA38);
	ND4 PPOO33(POO33, PAA39, PAA310, POO31, POO32);

	ND2 PPAA41(PAA41, Y04, Y14);
	ND2 PPAA42(PAA42, Y04, Y24);
	ND2 PPAA43(PAA43, Y04, Y34);
	ND2 PPAA44(PAA44, Y04, Y44);
	ND2 PPAA45(PAA45, Y14, Y24);
	ND2 PPAA46(PAA46, Y14, Y34);
	ND2 PPAA47(PAA47, Y14, Y44);
	ND2 PPAA48(PAA48, Y24, Y34);
	ND2 PPAA49(PAA49, Y24, Y44);
	ND2 PPAA410(PAA410, Y34, Y44);
	AN4 PPOO41(POO41, PAA41, PAA42, PAA43, PAA44);
	AN4 PPOO42(POO42, PAA45, PAA46, PAA47, PAA48);
	ND4 PPOO43(POO43, PAA49, PAA410, POO41, POO42);

	ND2 PPAA51(PAA51, Y05, Y15);
	ND2 PPAA52(PAA52, Y05, Y25);
	ND2 PPAA53(PAA53, Y05, Y35);
	ND2 PPAA54(PAA54, Y05, Y45);
	ND2 PPAA55(PAA55, Y15, Y25);
	ND2 PPAA56(PAA56, Y15, Y35);
	ND2 PPAA57(PAA57, Y15, Y45);
	ND2 PPAA58(PAA58, Y25, Y35);
	ND2 PPAA59(PAA59, Y25, Y45);
	ND2 PPAA510(PAA510, Y35, Y45);
	AN4 PPOO51(POO51, PAA51, PAA52, PAA53, PAA54);
	AN4 PPOO52(POO52, PAA55, PAA56, PAA57, PAA58);
	ND4 PPOO53(POO53, PAA59, PAA510, POO51, POO52);

	ND2 PPAA61(PAA61, Y06, Y16);
	ND2 PPAA62(PAA62, Y06, Y26);
	ND2 PPAA63(PAA63, Y06, Y36);
	ND2 PPAA64(PAA64, Y06, Y46);
	ND2 PPAA65(PAA65, Y16, Y26);
	ND2 PPAA66(PAA66, Y16, Y36);
	ND2 PPAA67(PAA67, Y16, Y46);
	ND2 PPAA68(PAA68, Y26, Y36);
	ND2 PPAA69(PAA69, Y26, Y46);
	ND2 PPAA610(PAA610, Y36, Y46);
	AN4 PPOO61(POO61, PAA61, PAA62, PAA63, PAA64);
	AN4 PPOO62(POO62, PAA65, PAA66, PAA67, PAA68);
	ND4 PPOO63(POO63, PAA69, PAA610, POO61, POO62);

	ND2 PPAA71(PAA71, Y07, Y17);
	ND2 PPAA72(PAA72, Y07, Y27);
	ND2 PPAA73(PAA73, Y07, Y37);
	ND2 PPAA74(PAA74, Y07, Y47);
	ND2 PPAA75(PAA75, Y17, Y27);
	ND2 PPAA76(PAA76, Y17, Y37);
	ND2 PPAA77(PAA77, Y17, Y47);
	ND2 PPAA78(PAA78, Y27, Y37);
	ND2 PPAA79(PAA79, Y27, Y47);
	ND2 PPAA710(PAA710, Y37, Y47);
	AN4 PPOO71(POO71, PAA71, PAA72, PAA73, PAA74);
	AN4 PPOO72(POO72, PAA75, PAA76, PAA77, PAA78);
	ND4 PPOO73(POO73, PAA79, PAA710, POO71, POO72);

	ND2 PPAA81(PAA81, Y08, Y18);
	ND2 PPAA82(PAA82, Y08, Y28);
	ND2 PPAA83(PAA83, Y08, Y38);
	ND2 PPAA84(PAA84, Y08, Y48);
	ND2 PPAA85(PAA85, Y18, Y28);
	ND2 PPAA86(PAA86, Y18, Y38);
	ND2 PPAA87(PAA87, Y18, Y48);
	ND2 PPAA88(PAA88, Y28, Y38);
	ND2 PPAA89(PAA89, Y28, Y48);
	ND2 PPAA810(PAA810, Y38, Y48);
	AN4 PPOO81(POO81, PAA81, PAA82, PAA83, PAA84);
	AN4 PPOO82(POO82, PAA85, PAA86, PAA87, PAA88);
	ND4 PPOO83(POO83, PAA89, PAA810, POO81, POO82);

	ND2 PPAA91(PAA91, Y09, Y19);
	ND2 PPAA92(PAA92, Y09, Y29);
	ND2 PPAA93(PAA93, Y09, Y39);
	ND2 PPAA94(PAA94, Y09, Y49);
	ND2 PPAA95(PAA95, Y19, Y29);
	ND2 PPAA96(PAA96, Y19, Y39);
	ND2 PPAA97(PAA97, Y19, Y49);
	ND2 PPAA98(PAA98, Y29, Y39);
	ND2 PPAA99(PAA99, Y29, Y49);
	ND2 PPAA910(PAA910, Y39, Y49);
	AN4 PPOO91(POO91, PAA91, PAA92, PAA93, PAA94);
	AN4 PPOO92(POO92, PAA95, PAA96, PAA97, PAA98);
	ND4 PPOO93(POO93, PAA99, PAA910, POO91, POO92);

	ND2 PPAA101(PAA101, Y010, Y110);
	ND2 PPAA102(PAA102, Y010, Y210);
	ND2 PPAA103(PAA103, Y010, Y310);
	ND2 PPAA104(PAA104, Y010, Y410);
	ND2 PPAA105(PAA105, Y110, Y210);
	ND2 PPAA106(PAA106, Y110, Y310);
	ND2 PPAA107(PAA107, Y110, Y410);
	ND2 PPAA108(PAA108, Y210, Y310);
	ND2 PPAA109(PAA109, Y210, Y410);
	ND2 PPAA1010(PAA1010, Y310, Y410);
	AN4 PPOO101(POO101, PAA101, PAA102, PAA103, PAA104);
	AN4 PPOO102(POO102, PAA105, PAA106, PAA107, PAA108);
	ND4 PPOO103(POO103, PAA109, PAA1010, POO101, POO102);

	ND2 PPAA111(PAA111, Y011, Y111);
	ND2 PPAA112(PAA112, Y011, Y211);
	ND2 PPAA113(PAA113, Y011, Y311);
	ND2 PPAA114(PAA114, Y011, Y411);
	ND2 PPAA115(PAA115, Y111, Y211);
	ND2 PPAA116(PAA116, Y111, Y311);
	ND2 PPAA117(PAA117, Y111, Y411);
	ND2 PPAA118(PAA118, Y211, Y311);
	ND2 PPAA119(PAA119, Y211, Y411);
	ND2 PPAA1110(PAA1110, Y311, Y411);
	AN4 PPOO111(POO111, PAA111, PAA112, PAA113, PAA114);
	AN4 PPOO112(POO112, PAA115, PAA116, PAA117, PAA118);
	ND4 PPOO113(POO113, PAA119, PAA1110, POO111, POO112);

	ND2 PPAA121(PAA121, Y012, Y112);
	ND2 PPAA122(PAA122, Y012, Y212);
	ND2 PPAA123(PAA123, Y012, Y312);
	ND2 PPAA124(PAA124, Y012, Y412);
	ND2 PPAA125(PAA125, Y112, Y212);
	ND2 PPAA126(PAA126, Y112, Y312);
	ND2 PPAA127(PAA127, Y112, Y412);
	ND2 PPAA128(PAA128, Y212, Y312);
	ND2 PPAA129(PAA129, Y212, Y412);
	ND2 PPAA1210(PAA1210, Y312, Y412);
	AN4 PPOO121(POO121, PAA121, PAA122, PAA123, PAA124);
	AN4 PPOO122(POO122, PAA125, PAA126, PAA127, PAA128);
	ND4 PPOO123(POO123, PAA129, PAA1210, POO121, POO122);

	ND2 PPAA131(PAA131, Y013, Y113);
	ND2 PPAA132(PAA132, Y013, Y213);
	ND2 PPAA133(PAA133, Y013, Y313);
	ND2 PPAA134(PAA134, Y013, Y413);
	ND2 PPAA135(PAA135, Y113, Y213);
	ND2 PPAA136(PAA136, Y113, Y313);
	ND2 PPAA137(PAA137, Y113, Y413);
	ND2 PPAA138(PAA138, Y213, Y313);
	ND2 PPAA139(PAA139, Y213, Y413);
	ND2 PPAA1310(PAA1310, Y313, Y413);
	AN4 PPOO131(POO131, PAA131, PAA132, PAA133, PAA134);
	AN4 PPOO132(POO132, PAA135, PAA136, PAA137, PAA138);
	ND4 PPOO133(POO133, PAA139, PAA1310, POO131, POO132);

	NR3 PPSS11(PSS11, POO13, POO23, POO33);
	NR3 PPSS21(PSS21, POO43, POO53, POO63);
	NR3 PPSS31(PSS31, POO73, POO83, POO93);
	NR4 PPSS41(PSS41, POO103, POO113, POO123, POO133);
	ND4 PPSS51(Q2, PSS11, PSS21, PSS31, PSS41);
	AN4 PPSS511(NQ2, PSS11, PSS21, PSS31, PSS41);

	ND4 PPAAA11(PAAA11, Y11, Y21, Y31, Y41);
	ND4 PPAAA12(PAAA12, Y01, Y21, Y31, Y41);
	ND4 PPAAA13(PAAA13, Y01, Y11, Y31, Y41);
	ND4 PPAAA14(PAAA14, Y01, Y11, Y21, Y41);
	ND4 PPAAA15(PAAA15, Y01, Y11, Y21, Y31);
	AN3 PPOOO11(POOO11, PAAA11, PAAA12, PAAA13);
	AN2 PPOOO12(POOO12, PAAA14, PAAA15);
	ND2 PPOOO13(POOO13, POOO11, POOO12);

	ND4 PPAAA21(PAAA21, Y12, Y22, Y32, Y42);
	ND4 PPAAA22(PAAA22, Y02, Y22, Y32, Y42);
	ND4 PPAAA23(PAAA23, Y02, Y12, Y32, Y42);
	ND4 PPAAA24(PAAA24, Y02, Y12, Y22, Y42);
	ND4 PPAAA25(PAAA25, Y02, Y12, Y22, Y32);
	AN3 PPOOO21(POOO21, PAAA21, PAAA22, PAAA23);
	AN2 PPOOO22(POOO22, PAAA24, PAAA25);
	ND2 PPOOO23(POOO23, POOO21, POOO22);

	ND4 PPAAA31(PAAA31, Y13, Y23, Y33, Y43);
	ND4 PPAAA32(PAAA32, Y03, Y23, Y33, Y43);
	ND4 PPAAA33(PAAA33, Y03, Y13, Y33, Y43);
	ND4 PPAAA34(PAAA34, Y03, Y13, Y23, Y43);
	ND4 PPAAA35(PAAA35, Y03, Y13, Y23, Y33);
	AN3 PPOOO31(POOO31, PAAA31, PAAA32, PAAA33);
	AN2 PPOOO32(POOO32, PAAA34, PAAA35);
	ND2 PPOOO33(POOO33, POOO31, POOO32);

	ND4 PPAAA41(PAAA41, Y14, Y24, Y34, Y44);
	ND4 PPAAA42(PAAA42, Y04, Y24, Y34, Y44);
	ND4 PPAAA43(PAAA43, Y04, Y14, Y34, Y44);
	ND4 PPAAA44(PAAA44, Y04, Y14, Y24, Y44);
	ND4 PPAAA45(PAAA45, Y04, Y14, Y24, Y34);
	AN3 PPOOO41(POOO41, PAAA41, PAAA42, PAAA43);
	AN2 PPOOO42(POOO42, PAAA44, PAAA45);
	ND2 PPOOO43(POOO43, POOO41, POOO42);

	ND4 PPAAA51(PAAA51, Y15, Y25, Y35, Y45);
	ND4 PPAAA52(PAAA52, Y05, Y25, Y35, Y45);
	ND4 PPAAA53(PAAA53, Y05, Y15, Y35, Y45);
	ND4 PPAAA54(PAAA54, Y05, Y15, Y25, Y45);
	ND4 PPAAA55(PAAA55, Y05, Y15, Y25, Y35);
	AN3 PPOOO51(POOO51, PAAA51, PAAA52, PAAA53);
	AN2 PPOOO52(POOO52, PAAA54, PAAA55);
	ND2 PPOOO53(POOO53, POOO51, POOO52);

	ND4 PPAAA61(PAAA61, Y16, Y26, Y36, Y46);
	ND4 PPAAA62(PAAA62, Y06, Y26, Y36, Y46);
	ND4 PPAAA63(PAAA63, Y06, Y16, Y36, Y46);
	ND4 PPAAA64(PAAA64, Y06, Y16, Y26, Y46);
	ND4 PPAAA65(PAAA65, Y06, Y16, Y26, Y36);
	AN3 PPOOO61(POOO61, PAAA61, PAAA62, PAAA63);
	AN2 PPOOO62(POOO62, PAAA64, PAAA65);
	ND2 PPOOO63(POOO63, POOO61, POOO62);

	ND4 PPAAA71(PAAA71, Y17, Y27, Y37, Y47);
	ND4 PPAAA72(PAAA72, Y07, Y27, Y37, Y47);
	ND4 PPAAA73(PAAA73, Y07, Y17, Y37, Y47);
	ND4 PPAAA74(PAAA74, Y07, Y17, Y27, Y47);
	ND4 PPAAA75(PAAA75, Y07, Y17, Y27, Y37);
	AN3 PPOOO71(POOO71, PAAA71, PAAA72, PAAA73);
	AN2 PPOOO72(POOO72, PAAA74, PAAA75);
	ND2 PPOOO73(POOO73, POOO71, POOO72);

	ND4 PPAAA81(PAAA81, Y18, Y28, Y38, Y48);
	ND4 PPAAA82(PAAA82, Y08, Y28, Y38, Y48);
	ND4 PPAAA83(PAAA83, Y08, Y18, Y38, Y48);
	ND4 PPAAA84(PAAA84, Y08, Y18, Y28, Y48);
	ND4 PPAAA85(PAAA85, Y08, Y18, Y28, Y38);
	AN3 PPOOO81(POOO81, PAAA81, PAAA82, PAAA83);
	AN2 PPOOO82(POOO82, PAAA84, PAAA85);
	ND2 PPOOO83(POOO83, POOO81, POOO82);

	ND4 PPAAA91(PAAA91, Y19, Y29, Y39, Y49);
	ND4 PPAAA92(PAAA92, Y09, Y29, Y39, Y49);
	ND4 PPAAA93(PAAA93, Y09, Y19, Y39, Y49);
	ND4 PPAAA94(PAAA94, Y09, Y19, Y29, Y49);
	ND4 PPAAA95(PAAA95, Y09, Y19, Y29, Y39);
	AN3 PPOOO91(POOO91, PAAA91, PAAA92, PAAA93);
	AN2 PPOOO92(POOO92, PAAA94, PAAA95);
	ND2 PPOOO93(POOO93, POOO91, POOO92);

	ND4 PPAAA101(PAAA101, Y110, Y210, Y310, Y410);
	ND4 PPAAA102(PAAA102, Y010, Y210, Y310, Y410);
	ND4 PPAAA103(PAAA103, Y010, Y110, Y310, Y410);
	ND4 PPAAA104(PAAA104, Y010, Y110, Y210, Y410);
	ND4 PPAAA105(PAAA105, Y010, Y110, Y210, Y310);
	AN3 PPOOO101(POOO101, PAAA101, PAAA102, PAAA103);
	AN2 PPOOO102(POOO102, PAAA104, PAAA105);
	ND2 PPOOO103(POOO103, POOO101, POOO102);

	ND4 PPAAA111(PAAA111, Y111, Y211, Y311, Y411);
	ND4 PPAAA112(PAAA112, Y011, Y211, Y311, Y411);
	ND4 PPAAA113(PAAA113, Y011, Y111, Y311, Y411);
	ND4 PPAAA114(PAAA114, Y011, Y111, Y211, Y411);
	ND4 PPAAA115(PAAA115, Y011, Y111, Y211, Y311);
	AN3 PPOOO111(POOO111, PAAA111, PAAA112, PAAA113);
	AN2 PPOOO112(POOO112, PAAA114, PAAA115);
	ND2 PPOOO113(POOO113, POOO111, POOO112);

	ND4 PPAAA121(PAAA121, Y112, Y212, Y312, Y412);
	ND4 PPAAA122(PAAA122, Y012, Y212, Y312, Y412);
	ND4 PPAAA123(PAAA123, Y012, Y112, Y312, Y412);
	ND4 PPAAA124(PAAA124, Y012, Y112, Y212, Y412);
	ND4 PPAAA125(PAAA125, Y012, Y112, Y212, Y312);
	AN3 PPOOO121(POOO121, PAAA121, PAAA122, PAAA123);
	AN2 PPOOO122(POOO122, PAAA124, PAAA125);
	ND2 PPOOO123(POOO123, POOO121, POOO122);

	ND4 PPAAA131(PAAA131, Y113, Y213, Y313, Y413);
	ND4 PPAAA132(PAAA132, Y013, Y213, Y313, Y413);
	ND4 PPAAA133(PAAA133, Y013, Y113, Y313, Y413);
	ND4 PPAAA134(PAAA134, Y013, Y113, Y213, Y413);
	ND4 PPAAA135(PAAA135, Y013, Y113, Y213, Y313);
	AN3 PPOOO131(POOO131, PAAA131, PAAA132, PAAA133);
	AN2 PPOOO132(POOO132, PAAA134, PAAA135);
	ND2 PPOOO133(POOO133, POOO131, POOO132);

	NR3 PPSSS11(PSSS11, POOO13, POOO23, POOO33);
	NR3 PPSSS21(PSSS21, POOO43, POOO53, POOO63);
	NR3 PPSSS31(PSSS31, POOO73, POOO83, POOO93);
	NR4 PPSSS41(PSSS41, POOO103, POOO113, POOO123, POOO133);
	ND4 PPSSS51(Q41, PSSS11, PSSS21, PSSS31, PSSS41);

	IV IVQ71(NPX71 ,PX71);
	IV L(NCHILL, CHILL);
	AN3 ANS32(Q32, Q3, Q2, NQ311);
	ND3 ANS322(NQ32, Q3, Q2, NQ311);
	AN3 ANS311(Q311, Q3, NQ221, PX71);
	ND3 ANS3111(NQ311, Q3, NQ221, PX71);
	AN3 ANS221(Q221, NPX71, NQ3, Q2);
	ND3 ANS2211(NQ221, NPX71, NQ3, Q2);
	AN3 ANS2111(Q2111, Q2, PX71, NQ3);
	AN2 ANS8(type[3], FLOWER, CHILL);
	AN2 ANS5(Q11111 , FLOWER, NCHILL);
	AN2 ANS4(J0, NF, CHILL);
	OR4 ANS2(type[2], Q11111, Q41, Q32, J0);
	OR4 ANS1(type[1], Q41, Q32, Q311, Q221);
	OR4 ANS0(type[0], Q41, Q311, Q2111, Q11111);

	EO3 PPX11(PX11, POO13, POO23, POO33);
	EO3 PPX21(PX21, POO43, POO53, POO63);
	EO3 PPX31(PX31, POO73, POO83, POO93);
	EO3 PPX41(PX41, POO103, POO113, POO123);
	EO3 PPX51(PX51, PX11, PX21, POO133);
	EO PPX61(PX61, PX31, PX41);
	EO PPX71(PX71, PX51, PX61);


endmodule